../../src/tlcWalk.vhd