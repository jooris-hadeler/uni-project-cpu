../../src/tlcTest.vhd