../../src/light.sv