src/de0Board.vhd