../../src/procPkg.vhd